library verilog;
use verilog.vl_types.all;
entity FixedPointAdder is
    port(
        in1             : in     vl_logic_vector(15 downto 0);
        in2             : in     vl_logic_vector(15 downto 0);
        \out\           : out    vl_logic_vector(15 downto 0)
    );
end FixedPointAdder;
