library verilog;
use verilog.vl_types.all;
entity TB_LDC is
end TB_LDC;
